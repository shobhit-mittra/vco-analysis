* CMOS-Inverter BAsed VCO - SPICE Netlist 

M1 N008 Fout N015 0 CMOSN l=180n w=540n
M2 N003 Fout N008 N001 CMOSP l=180n w=1350n
M3 N009 N008 N016 0 CMOSN l=180n w=540n
M4 N004 N008 N009 N001 CMOSP l=180n w=1350n
M5 N010 N009 N017 0 CMOSN l=180n w=540n
M6 N005 N009 N010 N001 CMOSP l=180n w=1350n
M7 N011 N010 N018 0 CMOSN l=180n w=540n
M8 N006 N010 N011 N001 CMOSP l=180n w=1350n
M9 Fout N011 N019 0 CMOSN l=180n w=540n
M10 N007 N011 Fout N001 CMOSP l=180n w=1350n
M11 N015 N020 0 0 CMOSN l=180n w=540n
M12 N016 N020 0 0 CMOSN l=180 w=540
M13 N017 N020 0 0 CMOSN l=180 w=540
M14 N018 N020 0 0 CMOSN l=180 w=540
M15 N019 N020 0 0 CMOSN l=180n w=540n
M16 N001 N002 N003 N001 CMOSP l=180n w=1350n
M17 N001 N002 N004 N001 CMOSP l=180n w=1350n
M18 N001 N002 N005 N001 CMOSP l=180n w=1350n
M19 N001 N002 N006 N001 CMOSP l=180n w=1350n
M20 N001 N002 N007 N001 CMOSP l=180n w=1350n
V1 N020 0 1
V2 N001 0 3
M21 N001 N002 N002 N001 CMOSP l=180n w=1350n
M22 N002 N020 0 0 CMOSN l=180n w=540n
M23 N012 Fout 0 0 CMOSN l=180n w=540n
M24 N001 Fout N012 N001 CMOSP l=180n w=1350n
M25 N013 N012 0 0 CMOSN l=180n w=540n
M26 N001 N012 N013 N001 CMOSP l=180n w=1350n
M27 N014 N013 0 0 CMOSN l=180n w=540n
M28 N001 N013 N014 N001 CMOSP l=180n w=1350n
M29 Fout_shaped N014 0 0 CMOSN l=180n w=540n
M30 N001 N014 Fout_shaped N001 CMOSP l=180n w=1350n
.model NMOS NMOS
.model PMOS PMOS
.lib ~\LTspiceXVII\lib\cmp\standard.mos  * Insert full path to standard mos lib on your system
.INCLUDE tsmc018.lib
* Diode Connected PMOS
* Vdd
* Vin
* Common Ground
.tran 15n
* Inverter stages for wave-shaping
.backanno
.end
